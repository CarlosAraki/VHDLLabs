--Nome:Carlos Vinícius Araki Oliveira RA:160141
--Nome:Cleber França Carvalho RA:145739

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EXP2a IS
	
	PORT ( SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
	
END EXP2a;

ARCHITECTURE Behavior OF EXP2a IS
	COMPONENT COMPARATOR IS
		PORT ( C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				  s: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT char_7seg
		PORT ( C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Display : OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	
	COMPONENT circA IS
	PORT ( C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			 S : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END COMPONENT;
	
COMPONENT circB IS
	PORT ( C : IN STD_LOGIC;
		 HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;

COMPONENT  Mux2_1 IS
	PORT ( x,y,s : IN STD_LOGIC;
			m : OUT STD_LOGIC);
	END COMPONENT ;

	SIGNAL Z,G,M0,M1,M2,M3: STD_LOGIC;
	SIGNAL VET: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL SEG: STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	BEGIN
	G <= '0';
	C0: COMPARATOR PORT MAP (SW(3 DOWNTO 0), Z);
	C1: circA PORT MAP (SW(2 DOWNTO 0), VET(2 DOWNTO 0));
	C2: mux2_1 PORT MAP(SW(0),VET(0),Z, M0);
	C3: mux2_1 PORT MAP(SW(1),VET(1),Z, M1);
	C4: mux2_1 PORT MAP(SW(2),VET(2),Z, M2);
	C5: mux2_1 PORT MAP(SW(3),G,Z, M3);
	C6: circB PORT MAP(Z,HEX1);
	SEG(0) <= M0;
	SEG(1) <= M1;
	SEG(2) <= M2;
	SEG(3) <= M3;
	C7: char_7seg PORT MAP(SEG,HEX0);
			
END Behavior;
