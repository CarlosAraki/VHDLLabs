--Nome:Carlos Vinícius Araki Oliveira RA:160141
--Nome:Cleber França Carvalho RA:145739

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EXP2a IS
	
	PORT ( SW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
	
END EXP2a;

ARCHITECTURE Behavior OF EXP2a IS


	COMPONENT COMPARATOR IS
	
	PORT ( C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 s: OUT STD_LOGIC);
	
	END COMPONENT;
	
	COMPONENT char_7seg
	PORT ( C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Display : OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	
	COMPONENT circA IS
	
	PORT ( C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			 S : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
	
END COMPONENT;
COMPONENT circB IS
	
	PORT ( C : IN STD_LOGIC;
			 HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
	
END COMPONENT;

	
	SIGNAL Z,M0,M1,M2,M3: STD_LOGIC;
		SIGNAL VECTORA: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL	VET1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	
	
	begin
	Q0 : COMPARATOR PORT MAP(SW(3 DOWNTO 0),Z);
	I0 : circA PORT MAP (SW(2 DOWNTO 0),VECTORA);
	M0 <= VECTORA(0) WHEN Z='1'
			ELSE SW(0);
	M1 <= VECTORA (1) WHEN Z='1'
			ELSE SW(1);
	M2 <= VECTORA (2) WHEN Z ='1'
			ELSE SW(2);
	M3 <= '0' WHEN Z='1'
			ELSE SW(3);
	VET1(0) <= M0;
	VET1(1) <= M1;
	VET1(2) <= M2;
	VET1(3) <= M3;
	O0:circB port map(Z,HEX1);
	P0: char_7seg PORT MAP(VET1,HEX0);
			
END Behavior;
